`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:24:11 02/01/2021 
// Design Name: 
// Module Name:    ActiveLamps 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ActiveLamps (
	input  [3:0] tcode        , // time code    [table2 time code   ]
	input  [3:0] ulight       , // user light   [light degree mode  ]
   input  [3:0] lenght       , // room length  [square room lenght ]
	output [3:0] active_lights  // number of active light
);

	reg [3:0] light_num;
	parameter morning = 4'b0001, afternoon = 4'b0010, evening = 4'b0100, night = 4'b1000;
	always @ (tcode or lenght or ulight)
		case(tcode)
			morning:   light_num =               4'b0000;
			afternoon: light_num =               4'b0000;
			evening:   light_num = {2'b00, lenght [3:2]}; // length*length/4*length = length/4
			night:     light_num =                ulight;
			default:   light_num =               4'b0000;
		endcase
	assign active_lights = light_num;
	
endmodule
